magic
tech sky130A
magscale 1 2
timestamp 1635942583
<< error_p >>
rect -2655 2230 -2429 2266
rect -2655 2148 -2619 2230
rect -2465 2148 -2429 2230
rect -2655 2112 -2429 2148
rect -1955 2230 -1729 2266
rect -1955 2148 -1919 2230
rect -1765 2148 -1729 2230
rect -1955 2112 -1729 2148
rect -1255 2230 -1029 2266
rect -1255 2148 -1219 2230
rect -1065 2148 -1029 2230
rect -1255 2112 -1029 2148
rect -555 2230 -329 2266
rect -555 2148 -519 2230
rect -365 2148 -329 2230
rect -555 2112 -329 2148
rect 145 2230 371 2266
rect 145 2148 181 2230
rect 335 2148 371 2230
rect 145 2112 371 2148
rect 845 2230 1071 2266
rect 845 2148 881 2230
rect 1035 2148 1071 2230
rect 845 2112 1071 2148
rect 1545 2230 1771 2266
rect 1545 2148 1581 2230
rect 1735 2148 1771 2230
rect 1545 2112 1771 2148
rect 2245 2230 2471 2266
rect 2245 2148 2281 2230
rect 2435 2148 2471 2230
rect 2245 2112 2471 2148
rect 2945 2230 3171 2266
rect 2945 2148 2981 2230
rect 3135 2148 3171 2230
rect 2945 2112 3171 2148
rect 3645 2230 3871 2266
rect 3645 2148 3681 2230
rect 3835 2148 3871 2230
rect 3645 2112 3871 2148
rect 5345 2230 5571 2266
rect 5345 2148 5381 2230
rect 5535 2148 5571 2230
rect 5345 2112 5571 2148
rect 6045 2230 6271 2266
rect 6045 2148 6081 2230
rect 6235 2148 6271 2230
rect 6045 2112 6271 2148
rect 6745 2230 6971 2266
rect 6745 2148 6781 2230
rect 6935 2148 6971 2230
rect 6745 2112 6971 2148
rect 7445 2230 7671 2266
rect 7445 2148 7481 2230
rect 7635 2148 7671 2230
rect 7445 2112 7671 2148
rect 8145 2230 8371 2266
rect 8145 2148 8181 2230
rect 8335 2148 8371 2230
rect 8145 2112 8371 2148
rect 8845 2230 9071 2266
rect 8845 2148 8881 2230
rect 9035 2148 9071 2230
rect 8845 2112 9071 2148
rect 9545 2230 9771 2266
rect 9545 2148 9581 2230
rect 9735 2148 9771 2230
rect 9545 2112 9771 2148
rect 10245 2230 10471 2266
rect 10245 2148 10281 2230
rect 10435 2148 10471 2230
rect 10245 2112 10471 2148
rect 10945 2230 11171 2266
rect 10945 2148 10981 2230
rect 11135 2148 11171 2230
rect 10945 2112 11171 2148
rect 11645 2230 11871 2266
rect 11645 2148 11681 2230
rect 11835 2148 11871 2230
rect 11645 2112 11871 2148
use m10_nfet_w10_l1  m10_nfet_w10_l1_0
array 0 1 8000 0 0 0
timestamp 1635942583
transform 1 0 -197 0 1 18
box -2712 -817 4234 2603
<< end >>
