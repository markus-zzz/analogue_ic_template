magic
tech sky130A
magscale 1 2
timestamp 1635942583
<< error_p >>
rect 15587 7010 15641 7144
rect 16335 7010 16541 7144
rect 17235 7010 17441 7144
rect 18135 7010 18341 7144
rect 14327 6383 14348 6915
rect 14384 6449 14414 6849
rect 14870 6449 14900 6849
rect 14936 6383 14966 6915
rect 15218 6383 15248 6915
rect 15284 6449 15314 6849
rect 15770 6449 15800 6849
rect 15836 6383 15866 6915
rect 16118 6383 16148 6915
rect 16184 6449 16214 6849
rect 16670 6449 16700 6849
rect 16736 6383 16766 6915
rect 17018 6383 17048 6915
rect 17084 6449 17114 6849
rect 17570 6449 17600 6849
rect 17636 6383 17666 6915
rect 17918 6383 17948 6915
rect 17984 6449 18014 6849
rect 18470 6449 18500 6849
rect 18536 6383 18566 6915
rect -4212 5949 -3986 5985
rect -4212 5867 -4176 5949
rect -4022 5867 -3986 5949
rect -4212 5831 -3986 5867
rect -3512 5949 -3286 5985
rect -3512 5867 -3476 5949
rect -3322 5867 -3286 5949
rect -3512 5831 -3286 5867
rect -2812 5949 -2586 5985
rect -2812 5867 -2776 5949
rect -2622 5867 -2586 5949
rect -2812 5831 -2586 5867
rect -2112 5949 -1886 5985
rect -2112 5867 -2076 5949
rect -1922 5867 -1886 5949
rect -2112 5831 -1886 5867
rect -1412 5949 -1346 5985
rect -1412 5867 -1376 5949
rect -1412 5831 -1346 5867
rect 14327 5643 14348 6175
rect 14384 5709 14414 6109
rect 14870 5709 14900 6109
rect 14936 5643 14966 6175
rect 15218 5643 15248 6175
rect 15284 5709 15314 6109
rect 15770 5709 15800 6109
rect 15836 5643 15866 6175
rect 16118 5643 16148 6175
rect 16184 5709 16214 6109
rect 16670 5709 16700 6109
rect 16736 5643 16766 6175
rect 17018 5643 17048 6175
rect 17084 5709 17114 6109
rect 17570 5709 17600 6109
rect 17636 5643 17666 6175
rect 17918 5643 17948 6175
rect 17984 5709 18014 6109
rect 18470 5709 18500 6109
rect 18536 5643 18566 6175
rect 15587 5405 15638 5539
rect 16332 5405 16538 5539
rect 17232 5405 17438 5539
rect 18132 5405 18338 5539
<< error_s >>
rect 2117 8670 2323 8804
rect 3117 8670 3323 8804
rect 1900 8043 1930 8575
rect 1966 8109 1996 8509
rect 2452 8109 2482 8509
rect 2518 8043 2548 8575
rect 2900 8043 2930 8575
rect 2966 8109 2996 8509
rect 3452 8109 3482 8509
rect 3518 8043 3548 8575
rect 1900 7303 1930 7835
rect 1966 7369 1996 7769
rect 2452 7369 2482 7769
rect 2518 7303 2548 7835
rect 2900 7303 2930 7835
rect 2966 7369 2996 7769
rect 3452 7369 3482 7769
rect 3518 7303 3548 7835
rect 2114 7065 2320 7199
rect 3114 7065 3320 7199
rect 11835 7010 12041 7144
rect 12735 7010 12941 7144
rect 13635 7010 13841 7144
rect 11618 6383 11648 6915
rect 11684 6449 11714 6849
rect 12170 6449 12200 6849
rect 12236 6383 12266 6915
rect 12518 6383 12548 6915
rect 12584 6449 12614 6849
rect 13070 6449 13100 6849
rect 13136 6383 13166 6915
rect 13418 6383 13448 6915
rect 13484 6449 13514 6849
rect 13970 6449 14000 6849
rect 14036 6383 14066 6915
rect 14318 6383 14327 6915
rect -1346 5949 -1186 5985
rect -1222 5867 -1186 5949
rect -1346 5831 -1186 5867
rect -712 5949 -486 5985
rect -712 5867 -676 5949
rect -522 5867 -486 5949
rect -712 5831 -486 5867
rect -12 5949 214 5985
rect -12 5867 24 5949
rect 178 5867 214 5949
rect -12 5831 214 5867
rect 688 5949 914 5985
rect 688 5867 724 5949
rect 878 5867 914 5949
rect 688 5831 914 5867
rect 1388 5949 1614 5985
rect 1388 5867 1424 5949
rect 1578 5867 1614 5949
rect 1388 5831 1614 5867
rect 2088 5949 2314 5985
rect 2088 5867 2124 5949
rect 2278 5867 2314 5949
rect 2088 5831 2314 5867
rect 3788 5949 4014 5985
rect 3788 5867 3824 5949
rect 3978 5867 4014 5949
rect 3788 5831 4014 5867
rect 4488 5949 4714 5985
rect 4488 5867 4524 5949
rect 4678 5867 4714 5949
rect 4488 5831 4714 5867
rect 5188 5949 5414 5985
rect 5188 5867 5224 5949
rect 5378 5867 5414 5949
rect 5188 5831 5414 5867
rect 5888 5949 6114 5985
rect 5888 5867 5924 5949
rect 6078 5867 6114 5949
rect 5888 5831 6114 5867
rect 6588 5949 6814 5985
rect 6588 5867 6624 5949
rect 6778 5867 6814 5949
rect 6588 5831 6814 5867
rect 7288 5949 7514 5985
rect 7288 5867 7324 5949
rect 7478 5867 7514 5949
rect 7288 5831 7514 5867
rect 7988 5949 8214 5985
rect 7988 5867 8024 5949
rect 8178 5867 8214 5949
rect 7988 5831 8214 5867
rect 8688 5949 8914 5985
rect 8688 5867 8724 5949
rect 8878 5867 8914 5949
rect 8688 5831 8914 5867
rect 9388 5949 9614 5985
rect 9388 5867 9424 5949
rect 9578 5867 9614 5949
rect 9388 5831 9614 5867
rect 10088 5949 10314 5985
rect 10088 5867 10124 5949
rect 10278 5867 10314 5949
rect 10088 5831 10314 5867
rect 11618 5643 11648 6175
rect 11684 5709 11714 6109
rect 12170 5709 12200 6109
rect 12236 5643 12266 6175
rect 12518 5643 12548 6175
rect 12584 5709 12614 6109
rect 13070 5709 13100 6109
rect 13136 5643 13166 6175
rect 13418 5643 13448 6175
rect 13484 5709 13514 6109
rect 13970 5709 14000 6109
rect 14036 5643 14066 6175
rect 14318 5643 14327 6175
rect 11832 5405 12038 5539
rect 12732 5405 12938 5539
rect 13632 5405 13838 5539
rect 1225 2158 1451 2194
rect 1225 2076 1261 2158
rect 1415 2076 1451 2158
rect 1225 2040 1451 2076
rect 2225 2158 2451 2194
rect 2225 2076 2261 2158
rect 2415 2076 2451 2158
rect 2225 2040 2451 2076
rect 3225 2158 3451 2194
rect 3225 2076 3261 2158
rect 3415 2076 3451 2158
rect 3225 2040 3451 2076
rect 4225 2158 4451 2194
rect 4225 2076 4261 2158
rect 4415 2076 4451 2158
rect 4225 2040 4451 2076
rect 5225 2158 5451 2194
rect 5225 2076 5261 2158
rect 5415 2076 5451 2158
rect 5225 2040 5451 2076
rect 6225 2158 6451 2194
rect 6225 2076 6261 2158
rect 6415 2076 6451 2158
rect 6225 2040 6451 2076
rect 7225 2158 7451 2194
rect 7225 2076 7261 2158
rect 7415 2076 7451 2158
rect 7225 2040 7451 2076
rect 8225 2158 8451 2194
rect 8225 2076 8261 2158
rect 8415 2076 8451 2158
rect 8225 2040 8451 2076
rect 9225 2158 9451 2194
rect 9225 2076 9261 2158
rect 9415 2076 9451 2158
rect 9225 2040 9451 2076
rect 10225 2158 10451 2194
rect 10225 2076 10261 2158
rect 10415 2076 10451 2158
rect 10225 2040 10451 2076
rect 1224 1021 1450 1057
rect 1224 939 1260 1021
rect 1414 939 1450 1021
rect 1224 903 1450 939
rect 2224 1021 2450 1057
rect 2224 939 2260 1021
rect 2414 939 2450 1021
rect 2224 903 2450 939
rect 3224 1021 3450 1057
rect 3224 939 3260 1021
rect 3414 939 3450 1021
rect 3224 903 3450 939
rect 4224 1021 4450 1057
rect 4224 939 4260 1021
rect 4414 939 4450 1021
rect 4224 903 4450 939
rect 5224 1021 5450 1057
rect 5224 939 5260 1021
rect 5414 939 5450 1021
rect 5224 903 5450 939
rect 6224 1021 6450 1057
rect 6224 939 6260 1021
rect 6414 939 6450 1021
rect 6224 903 6450 939
rect 7224 1021 7450 1057
rect 7224 939 7260 1021
rect 7414 939 7450 1021
rect 7224 903 7450 939
rect 8224 1021 8450 1057
rect 8224 939 8260 1021
rect 8414 939 8450 1021
rect 8224 903 8450 939
rect 9224 1021 9450 1057
rect 9224 939 9260 1021
rect 9414 939 9450 1021
rect 9224 903 9450 939
rect 10224 1021 10450 1057
rect 10224 939 10260 1021
rect 10414 939 10450 1021
rect 10224 903 10450 939
<< error_ps >>
rect 14535 7010 14741 7144
rect 15435 7010 15587 7144
rect 14532 5405 14738 5539
rect 15432 5405 15587 5539
<< metal1 >>
rect 1551 8950 1669 9069
rect 2972 8951 4266 9070
rect 4125 7474 4266 8951
rect 4125 7291 11226 7474
rect 2476 6413 2609 6910
rect 2012 6182 2614 6413
rect 3476 6409 3609 6910
rect 3477 6188 3609 6409
rect 12291 3975 12461 5064
rect 12291 3621 13067 3975
rect 2480 2920 4044 3080
rect 956 2287 1083 2411
rect 2586 2397 2711 2920
rect 12291 2520 12461 3621
rect 10711 2397 12461 2520
rect 652 495 852 713
<< metal2 >>
rect 9880 6229 11838 6329
rect -86 5849 60 5951
rect 3845 5849 3991 5951
rect 1786 3404 1937 3492
rect 9752 3405 9920 3493
use contact$4  contact$4_0
timestamp 1635942583
transform 1 0 9996 0 1 6278
box -64 -32 64 32
use diff_pair  diff_pair_0
timestamp 1635942583
transform 1 0 -1557 0 1 3719
box -2909 -799 12037 2621
use current_mirror  current_mirror_0
timestamp 1635942583
transform 1 0 2847 0 1 7379
box -1298 -469 762 1691
use amp  amp_0
timestamp 1635942583
transform 1 0 14597 0 1 6161
box -3371 -1097 4030 1313
use bias_current_mirror  bias_current_mirror_0
timestamp 1635942583
transform 1 0 2122 0 1 3452
box -1470 -2957 8696 488
<< labels >>
flabel metal1 s 1551 8950 1669 9069 2 FreeSans 2000 0 0 0 vdd
port 1 nsew
flabel metal1 s 12747 3625 13063 3972 2 FreeSans 2000 0 0 0 out
port 2 nsew
flabel metal1 s 652 495 852 713 2 FreeSans 2000 0 0 0 vss
port 3 nsew
flabel metal1 s 956 2287 1083 2411 2 FreeSans 2000 0 0 0 bias
port 4 nsew
flabel metal2 s 1786 3404 1937 3492 2 FreeSans 2000 0 0 0 in_n
port 5 nsew
flabel metal2 s 9752 3405 9920 3493 2 FreeSans 2000 0 0 0 in_p
port 6 nsew
flabel metal2 s 3845 5849 3991 5951 2 FreeSans 2000 0 0 0 vss
port 3 nsew
flabel metal2 s -86 5849 60 5951 2 FreeSans 2000 0 0 0 vss
port 3 nsew
<< end >>
