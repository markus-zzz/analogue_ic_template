magic
tech sky130A
magscale 1 2
timestamp 1635942583
<< error_s >>
rect -107 1101 99 1235
rect -324 474 -294 1006
rect -258 540 -228 940
rect 228 540 258 940
rect 294 474 324 1006
rect -324 -266 -294 266
rect -258 -200 -228 200
rect 228 -200 258 200
rect 294 -266 324 266
rect -110 -504 96 -370
<< metal1 >>
rect -385 1220 -252 1382
rect -385 1116 76 1220
rect -385 -385 -252 1116
rect -196 287 196 453
rect -385 -489 76 -385
rect 252 -659 385 1071
use sky130_fd_pr__pfet_g5v0d10v5_QSRSHK  sky130_fd_pr__pfet_g5v0d10v5_QSRSHK_0
array 0 0 0 0 1 740
timestamp 1635942583
transform 1 0 0 0 1 0
box -324 -576 324 534
use contact$3  contact$3_0
timestamp 1635942583
transform 1 0 -4 0 1 1168
box -69 -33 69 33
use contact$2  contact$2_0
timestamp 1635942583
transform 1 0 -4 0 1 1168
box -103 -67 103 67
use contact$3  contact$3_1
timestamp 1635942583
transform 1 0 -7 0 1 -437
box -69 -33 69 33
use contact$2  contact$2_1
timestamp 1635942583
transform 1 0 -7 0 1 -437
box -103 -67 103 67
<< end >>
