magic
tech sky130A
magscale 1 2
timestamp 1635942583
<< pwell >>
rect -184 -1026 184 1026
<< mvnmos >>
rect -100 -1000 100 1000
<< mvndiff >>
rect -158 969 -100 1000
rect -158 935 -146 969
rect -112 935 -100 969
rect -158 901 -100 935
rect -158 867 -146 901
rect -112 867 -100 901
rect -158 833 -100 867
rect -158 799 -146 833
rect -112 799 -100 833
rect -158 765 -100 799
rect -158 731 -146 765
rect -112 731 -100 765
rect -158 697 -100 731
rect -158 663 -146 697
rect -112 663 -100 697
rect -158 629 -100 663
rect -158 595 -146 629
rect -112 595 -100 629
rect -158 561 -100 595
rect -158 527 -146 561
rect -112 527 -100 561
rect -158 493 -100 527
rect -158 459 -146 493
rect -112 459 -100 493
rect -158 425 -100 459
rect -158 391 -146 425
rect -112 391 -100 425
rect -158 357 -100 391
rect -158 323 -146 357
rect -112 323 -100 357
rect -158 289 -100 323
rect -158 255 -146 289
rect -112 255 -100 289
rect -158 221 -100 255
rect -158 187 -146 221
rect -112 187 -100 221
rect -158 153 -100 187
rect -158 119 -146 153
rect -112 119 -100 153
rect -158 85 -100 119
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -119 -100 -85
rect -158 -153 -146 -119
rect -112 -153 -100 -119
rect -158 -187 -100 -153
rect -158 -221 -146 -187
rect -112 -221 -100 -187
rect -158 -255 -100 -221
rect -158 -289 -146 -255
rect -112 -289 -100 -255
rect -158 -323 -100 -289
rect -158 -357 -146 -323
rect -112 -357 -100 -323
rect -158 -391 -100 -357
rect -158 -425 -146 -391
rect -112 -425 -100 -391
rect -158 -459 -100 -425
rect -158 -493 -146 -459
rect -112 -493 -100 -459
rect -158 -527 -100 -493
rect -158 -561 -146 -527
rect -112 -561 -100 -527
rect -158 -595 -100 -561
rect -158 -629 -146 -595
rect -112 -629 -100 -595
rect -158 -663 -100 -629
rect -158 -697 -146 -663
rect -112 -697 -100 -663
rect -158 -731 -100 -697
rect -158 -765 -146 -731
rect -112 -765 -100 -731
rect -158 -799 -100 -765
rect -158 -833 -146 -799
rect -112 -833 -100 -799
rect -158 -867 -100 -833
rect -158 -901 -146 -867
rect -112 -901 -100 -867
rect -158 -935 -100 -901
rect -158 -969 -146 -935
rect -112 -969 -100 -935
rect -158 -1000 -100 -969
rect 100 969 158 1000
rect 100 935 112 969
rect 146 935 158 969
rect 100 901 158 935
rect 100 867 112 901
rect 146 867 158 901
rect 100 833 158 867
rect 100 799 112 833
rect 146 799 158 833
rect 100 765 158 799
rect 100 731 112 765
rect 146 731 158 765
rect 100 697 158 731
rect 100 663 112 697
rect 146 663 158 697
rect 100 629 158 663
rect 100 595 112 629
rect 146 595 158 629
rect 100 561 158 595
rect 100 527 112 561
rect 146 527 158 561
rect 100 493 158 527
rect 100 459 112 493
rect 146 459 158 493
rect 100 425 158 459
rect 100 391 112 425
rect 146 391 158 425
rect 100 357 158 391
rect 100 323 112 357
rect 146 323 158 357
rect 100 289 158 323
rect 100 255 112 289
rect 146 255 158 289
rect 100 221 158 255
rect 100 187 112 221
rect 146 187 158 221
rect 100 153 158 187
rect 100 119 112 153
rect 146 119 158 153
rect 100 85 158 119
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -119 158 -85
rect 100 -153 112 -119
rect 146 -153 158 -119
rect 100 -187 158 -153
rect 100 -221 112 -187
rect 146 -221 158 -187
rect 100 -255 158 -221
rect 100 -289 112 -255
rect 146 -289 158 -255
rect 100 -323 158 -289
rect 100 -357 112 -323
rect 146 -357 158 -323
rect 100 -391 158 -357
rect 100 -425 112 -391
rect 146 -425 158 -391
rect 100 -459 158 -425
rect 100 -493 112 -459
rect 146 -493 158 -459
rect 100 -527 158 -493
rect 100 -561 112 -527
rect 146 -561 158 -527
rect 100 -595 158 -561
rect 100 -629 112 -595
rect 146 -629 158 -595
rect 100 -663 158 -629
rect 100 -697 112 -663
rect 146 -697 158 -663
rect 100 -731 158 -697
rect 100 -765 112 -731
rect 146 -765 158 -731
rect 100 -799 158 -765
rect 100 -833 112 -799
rect 146 -833 158 -799
rect 100 -867 158 -833
rect 100 -901 112 -867
rect 146 -901 158 -867
rect 100 -935 158 -901
rect 100 -969 112 -935
rect 146 -969 158 -935
rect 100 -1000 158 -969
<< mvndiffc >>
rect -146 935 -112 969
rect -146 867 -112 901
rect -146 799 -112 833
rect -146 731 -112 765
rect -146 663 -112 697
rect -146 595 -112 629
rect -146 527 -112 561
rect -146 459 -112 493
rect -146 391 -112 425
rect -146 323 -112 357
rect -146 255 -112 289
rect -146 187 -112 221
rect -146 119 -112 153
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect -146 -153 -112 -119
rect -146 -221 -112 -187
rect -146 -289 -112 -255
rect -146 -357 -112 -323
rect -146 -425 -112 -391
rect -146 -493 -112 -459
rect -146 -561 -112 -527
rect -146 -629 -112 -595
rect -146 -697 -112 -663
rect -146 -765 -112 -731
rect -146 -833 -112 -799
rect -146 -901 -112 -867
rect -146 -969 -112 -935
rect 112 935 146 969
rect 112 867 146 901
rect 112 799 146 833
rect 112 731 146 765
rect 112 663 146 697
rect 112 595 146 629
rect 112 527 146 561
rect 112 459 146 493
rect 112 391 146 425
rect 112 323 146 357
rect 112 255 146 289
rect 112 187 146 221
rect 112 119 146 153
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
rect 112 -153 146 -119
rect 112 -221 146 -187
rect 112 -289 146 -255
rect 112 -357 146 -323
rect 112 -425 146 -391
rect 112 -493 146 -459
rect 112 -561 146 -527
rect 112 -629 146 -595
rect 112 -697 146 -663
rect 112 -765 146 -731
rect 112 -833 146 -799
rect 112 -901 146 -867
rect 112 -969 146 -935
<< poly >>
rect -100 1072 100 1088
rect -100 1038 -51 1072
rect -17 1038 17 1072
rect 51 1038 100 1072
rect -100 1000 100 1038
rect -100 -1038 100 -1000
rect -100 -1072 -51 -1038
rect -17 -1072 17 -1038
rect 51 -1072 100 -1038
rect -100 -1088 100 -1072
<< polycont >>
rect -51 1038 -17 1072
rect 17 1038 51 1072
rect -51 -1072 -17 -1038
rect 17 -1072 51 -1038
<< locali >>
rect -100 1038 -53 1072
rect -17 1038 17 1072
rect 53 1038 100 1072
rect -146 969 -112 1004
rect -146 901 -112 919
rect -146 833 -112 847
rect -146 765 -112 775
rect -146 697 -112 703
rect -146 629 -112 631
rect -146 593 -112 595
rect -146 521 -112 527
rect -146 449 -112 459
rect -146 377 -112 391
rect -146 305 -112 323
rect -146 233 -112 255
rect -146 161 -112 187
rect -146 89 -112 119
rect -146 17 -112 51
rect -146 -51 -112 -17
rect -146 -119 -112 -89
rect -146 -187 -112 -161
rect -146 -255 -112 -233
rect -146 -323 -112 -305
rect -146 -391 -112 -377
rect -146 -459 -112 -449
rect -146 -527 -112 -521
rect -146 -595 -112 -593
rect -146 -631 -112 -629
rect -146 -703 -112 -697
rect -146 -775 -112 -765
rect -146 -847 -112 -833
rect -146 -919 -112 -901
rect -146 -1004 -112 -969
rect 112 969 146 1004
rect 112 901 146 919
rect 112 833 146 847
rect 112 765 146 775
rect 112 697 146 703
rect 112 629 146 631
rect 112 593 146 595
rect 112 521 146 527
rect 112 449 146 459
rect 112 377 146 391
rect 112 305 146 323
rect 112 233 146 255
rect 112 161 146 187
rect 112 89 146 119
rect 112 17 146 51
rect 112 -51 146 -17
rect 112 -119 146 -89
rect 112 -187 146 -161
rect 112 -255 146 -233
rect 112 -323 146 -305
rect 112 -391 146 -377
rect 112 -459 146 -449
rect 112 -527 146 -521
rect 112 -595 146 -593
rect 112 -631 146 -629
rect 112 -703 146 -697
rect 112 -775 146 -765
rect 112 -847 146 -833
rect 112 -919 146 -901
rect 112 -1004 146 -969
rect -100 -1072 -53 -1038
rect -17 -1072 17 -1038
rect 53 -1072 100 -1038
<< viali >>
rect -53 1038 -51 1072
rect -51 1038 -19 1072
rect 19 1038 51 1072
rect 51 1038 53 1072
rect -146 935 -112 953
rect -146 919 -112 935
rect -146 867 -112 881
rect -146 847 -112 867
rect -146 799 -112 809
rect -146 775 -112 799
rect -146 731 -112 737
rect -146 703 -112 731
rect -146 663 -112 665
rect -146 631 -112 663
rect -146 561 -112 593
rect -146 559 -112 561
rect -146 493 -112 521
rect -146 487 -112 493
rect -146 425 -112 449
rect -146 415 -112 425
rect -146 357 -112 377
rect -146 343 -112 357
rect -146 289 -112 305
rect -146 271 -112 289
rect -146 221 -112 233
rect -146 199 -112 221
rect -146 153 -112 161
rect -146 127 -112 153
rect -146 85 -112 89
rect -146 55 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -55
rect -146 -89 -112 -85
rect -146 -153 -112 -127
rect -146 -161 -112 -153
rect -146 -221 -112 -199
rect -146 -233 -112 -221
rect -146 -289 -112 -271
rect -146 -305 -112 -289
rect -146 -357 -112 -343
rect -146 -377 -112 -357
rect -146 -425 -112 -415
rect -146 -449 -112 -425
rect -146 -493 -112 -487
rect -146 -521 -112 -493
rect -146 -561 -112 -559
rect -146 -593 -112 -561
rect -146 -663 -112 -631
rect -146 -665 -112 -663
rect -146 -731 -112 -703
rect -146 -737 -112 -731
rect -146 -799 -112 -775
rect -146 -809 -112 -799
rect -146 -867 -112 -847
rect -146 -881 -112 -867
rect -146 -935 -112 -919
rect -146 -953 -112 -935
rect 112 935 146 953
rect 112 919 146 935
rect 112 867 146 881
rect 112 847 146 867
rect 112 799 146 809
rect 112 775 146 799
rect 112 731 146 737
rect 112 703 146 731
rect 112 663 146 665
rect 112 631 146 663
rect 112 561 146 593
rect 112 559 146 561
rect 112 493 146 521
rect 112 487 146 493
rect 112 425 146 449
rect 112 415 146 425
rect 112 357 146 377
rect 112 343 146 357
rect 112 289 146 305
rect 112 271 146 289
rect 112 221 146 233
rect 112 199 146 221
rect 112 153 146 161
rect 112 127 146 153
rect 112 85 146 89
rect 112 55 146 85
rect 112 -17 146 17
rect 112 -85 146 -55
rect 112 -89 146 -85
rect 112 -153 146 -127
rect 112 -161 146 -153
rect 112 -221 146 -199
rect 112 -233 146 -221
rect 112 -289 146 -271
rect 112 -305 146 -289
rect 112 -357 146 -343
rect 112 -377 146 -357
rect 112 -425 146 -415
rect 112 -449 146 -425
rect 112 -493 146 -487
rect 112 -521 146 -493
rect 112 -561 146 -559
rect 112 -593 146 -561
rect 112 -663 146 -631
rect 112 -665 146 -663
rect 112 -731 146 -703
rect 112 -737 146 -731
rect 112 -799 146 -775
rect 112 -809 146 -799
rect 112 -867 146 -847
rect 112 -881 146 -867
rect 112 -935 146 -919
rect 112 -953 146 -935
rect -53 -1072 -51 -1038
rect -51 -1072 -19 -1038
rect 19 -1072 51 -1038
rect 51 -1072 53 -1038
<< metal1 >>
rect -96 1072 96 1078
rect -96 1038 -53 1072
rect -19 1038 19 1072
rect 53 1038 96 1072
rect -96 1032 96 1038
rect -152 953 -106 1000
rect -152 919 -146 953
rect -112 919 -106 953
rect -152 881 -106 919
rect -152 847 -146 881
rect -112 847 -106 881
rect -152 809 -106 847
rect -152 775 -146 809
rect -112 775 -106 809
rect -152 737 -106 775
rect -152 703 -146 737
rect -112 703 -106 737
rect -152 665 -106 703
rect -152 631 -146 665
rect -112 631 -106 665
rect -152 593 -106 631
rect -152 559 -146 593
rect -112 559 -106 593
rect -152 521 -106 559
rect -152 487 -146 521
rect -112 487 -106 521
rect -152 449 -106 487
rect -152 415 -146 449
rect -112 415 -106 449
rect -152 377 -106 415
rect -152 343 -146 377
rect -112 343 -106 377
rect -152 305 -106 343
rect -152 271 -146 305
rect -112 271 -106 305
rect -152 233 -106 271
rect -152 199 -146 233
rect -112 199 -106 233
rect -152 161 -106 199
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -199 -106 -161
rect -152 -233 -146 -199
rect -112 -233 -106 -199
rect -152 -271 -106 -233
rect -152 -305 -146 -271
rect -112 -305 -106 -271
rect -152 -343 -106 -305
rect -152 -377 -146 -343
rect -112 -377 -106 -343
rect -152 -415 -106 -377
rect -152 -449 -146 -415
rect -112 -449 -106 -415
rect -152 -487 -106 -449
rect -152 -521 -146 -487
rect -112 -521 -106 -487
rect -152 -559 -106 -521
rect -152 -593 -146 -559
rect -112 -593 -106 -559
rect -152 -631 -106 -593
rect -152 -665 -146 -631
rect -112 -665 -106 -631
rect -152 -703 -106 -665
rect -152 -737 -146 -703
rect -112 -737 -106 -703
rect -152 -775 -106 -737
rect -152 -809 -146 -775
rect -112 -809 -106 -775
rect -152 -847 -106 -809
rect -152 -881 -146 -847
rect -112 -881 -106 -847
rect -152 -919 -106 -881
rect -152 -953 -146 -919
rect -112 -953 -106 -919
rect -152 -1000 -106 -953
rect 106 953 152 1000
rect 106 919 112 953
rect 146 919 152 953
rect 106 881 152 919
rect 106 847 112 881
rect 146 847 152 881
rect 106 809 152 847
rect 106 775 112 809
rect 146 775 152 809
rect 106 737 152 775
rect 106 703 112 737
rect 146 703 152 737
rect 106 665 152 703
rect 106 631 112 665
rect 146 631 152 665
rect 106 593 152 631
rect 106 559 112 593
rect 146 559 152 593
rect 106 521 152 559
rect 106 487 112 521
rect 146 487 152 521
rect 106 449 152 487
rect 106 415 112 449
rect 146 415 152 449
rect 106 377 152 415
rect 106 343 112 377
rect 146 343 152 377
rect 106 305 152 343
rect 106 271 112 305
rect 146 271 152 305
rect 106 233 152 271
rect 106 199 112 233
rect 146 199 152 233
rect 106 161 152 199
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -199 152 -161
rect 106 -233 112 -199
rect 146 -233 152 -199
rect 106 -271 152 -233
rect 106 -305 112 -271
rect 146 -305 152 -271
rect 106 -343 152 -305
rect 106 -377 112 -343
rect 146 -377 152 -343
rect 106 -415 152 -377
rect 106 -449 112 -415
rect 146 -449 152 -415
rect 106 -487 152 -449
rect 106 -521 112 -487
rect 146 -521 152 -487
rect 106 -559 152 -521
rect 106 -593 112 -559
rect 146 -593 152 -559
rect 106 -631 152 -593
rect 106 -665 112 -631
rect 146 -665 152 -631
rect 106 -703 152 -665
rect 106 -737 112 -703
rect 146 -737 152 -703
rect 106 -775 152 -737
rect 106 -809 112 -775
rect 146 -809 152 -775
rect 106 -847 152 -809
rect 106 -881 112 -847
rect 146 -881 152 -847
rect 106 -919 152 -881
rect 106 -953 112 -919
rect 146 -953 152 -919
rect 106 -1000 152 -953
rect -96 -1038 96 -1032
rect -96 -1072 -53 -1038
rect -19 -1072 19 -1038
rect 53 -1072 96 -1038
rect -96 -1078 96 -1072
<< end >>
