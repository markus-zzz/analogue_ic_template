magic
tech sky130A
timestamp 1635942583
<< end >>
