magic
tech sky130A
magscale 1 2
timestamp 1635942583
<< error_s >>
rect -2458 2212 -2232 2248
rect -2458 2130 -2422 2212
rect -2268 2130 -2232 2212
rect -2458 2094 -2232 2130
rect -1758 2212 -1532 2248
rect -1758 2130 -1722 2212
rect -1568 2130 -1532 2212
rect -1758 2094 -1532 2130
rect -1058 2212 -832 2248
rect -1058 2130 -1022 2212
rect -868 2130 -832 2212
rect -1058 2094 -832 2130
rect -358 2212 -132 2248
rect -358 2130 -322 2212
rect -168 2130 -132 2212
rect -358 2094 -132 2130
rect 342 2212 568 2248
rect 342 2130 378 2212
rect 532 2130 568 2212
rect 342 2094 568 2130
rect 1042 2212 1268 2248
rect 1042 2130 1078 2212
rect 1232 2130 1268 2212
rect 1042 2094 1268 2130
rect 1742 2212 1968 2248
rect 1742 2130 1778 2212
rect 1932 2130 1968 2212
rect 1742 2094 1968 2130
rect 2442 2212 2668 2248
rect 2442 2130 2478 2212
rect 2632 2130 2668 2212
rect 2442 2094 2668 2130
rect 3142 2212 3368 2248
rect 3142 2130 3178 2212
rect 3332 2130 3368 2212
rect 3142 2094 3368 2130
rect 3842 2212 4068 2248
rect 3842 2130 3878 2212
rect 4032 2130 4068 2212
rect 3842 2094 4068 2130
<< metal1 >>
rect -2642 2443 3794 2603
rect -2202 -817 4234 -657
<< metal2 >>
rect -2712 2116 4043 2216
rect -2427 -323 4027 -238
use nfet_w10_l1  nfet_w10_l1_0
array 0 9 700 0 0 0
timestamp 1635942583
transform 1 0 372 0 1 99
box -3014 -756 -2438 2344
<< end >>
