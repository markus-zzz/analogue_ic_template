magic
tech sky130A
magscale 1 2
timestamp 1635942583
<< error_s >>
rect -897 -1294 -671 -1258
rect -897 -1376 -861 -1294
rect -707 -1376 -671 -1294
rect -897 -1412 -671 -1376
rect 103 -1294 329 -1258
rect 103 -1376 139 -1294
rect 293 -1376 329 -1294
rect 103 -1412 329 -1376
rect 1103 -1294 1329 -1258
rect 1103 -1376 1139 -1294
rect 1293 -1376 1329 -1294
rect 1103 -1412 1329 -1376
rect 2103 -1294 2329 -1258
rect 2103 -1376 2139 -1294
rect 2293 -1376 2329 -1294
rect 2103 -1412 2329 -1376
rect 3103 -1294 3329 -1258
rect 3103 -1376 3139 -1294
rect 3293 -1376 3329 -1294
rect 3103 -1412 3329 -1376
rect 4103 -1294 4329 -1258
rect 4103 -1376 4139 -1294
rect 4293 -1376 4329 -1294
rect 4103 -1412 4329 -1376
rect 5103 -1294 5329 -1258
rect 5103 -1376 5139 -1294
rect 5293 -1376 5329 -1294
rect 5103 -1412 5329 -1376
rect 6103 -1294 6329 -1258
rect 6103 -1376 6139 -1294
rect 6293 -1376 6329 -1294
rect 6103 -1412 6329 -1376
rect 7103 -1294 7329 -1258
rect 7103 -1376 7139 -1294
rect 7293 -1376 7329 -1294
rect 7103 -1412 7329 -1376
rect 8103 -1294 8329 -1258
rect 8103 -1376 8139 -1294
rect 8293 -1376 8329 -1294
rect 8103 -1412 8329 -1376
rect -898 -2431 -672 -2395
rect -898 -2513 -862 -2431
rect -708 -2513 -672 -2431
rect -898 -2549 -672 -2513
rect 102 -2431 328 -2395
rect 102 -2513 138 -2431
rect 292 -2513 328 -2431
rect 102 -2549 328 -2513
rect 1102 -2431 1328 -2395
rect 1102 -2513 1138 -2431
rect 1292 -2513 1328 -2431
rect 1102 -2549 1328 -2513
rect 2102 -2431 2328 -2395
rect 2102 -2513 2138 -2431
rect 2292 -2513 2328 -2431
rect 2102 -2549 2328 -2513
rect 3102 -2431 3328 -2395
rect 3102 -2513 3138 -2431
rect 3292 -2513 3328 -2431
rect 3102 -2549 3328 -2513
rect 4102 -2431 4328 -2395
rect 4102 -2513 4138 -2431
rect 4292 -2513 4328 -2431
rect 4102 -2549 4328 -2513
rect 5102 -2431 5328 -2395
rect 5102 -2513 5138 -2431
rect 5292 -2513 5328 -2431
rect 5102 -2549 5328 -2513
rect 6102 -2431 6328 -2395
rect 6102 -2513 6138 -2431
rect 6292 -2513 6328 -2431
rect 6102 -2549 6328 -2513
rect 7102 -2431 7328 -2395
rect 7102 -2513 7138 -2431
rect 7292 -2513 7328 -2431
rect 7102 -2549 7328 -2513
rect 8102 -2431 8328 -2395
rect 8102 -2513 8138 -2431
rect 8292 -2513 8328 -2431
rect 8102 -2549 8328 -2513
<< metal1 >>
rect -1166 -1165 -411 -1041
rect 1464 -1055 8589 -932
rect -536 -1395 -411 -1165
rect 464 -1395 589 -1055
rect 1464 -1395 1589 -1055
rect 2464 -1395 2589 -1055
rect 3464 -1395 3589 -1055
rect 4464 -1395 4589 -1055
rect 5464 -1395 5589 -1055
rect 6464 -1395 6589 -1055
rect 7464 -1395 7589 -1055
rect 8464 -1395 8589 -1055
rect -592 -1959 -536 -1815
rect -1470 -2957 8696 -2739
<< metal2 >>
rect -854 -1927 8305 -1843
use contact  contact_0
timestamp 1635942583
transform 1 0 -548 0 1 487
box 0 0 1 1
use m2_nfet_w1_l2  m2_nfet_w1_l2_0
array 0 9 1000 0 0 0
timestamp 1635942583
transform 1 0 -514 0 1 -1928
box -651 -811 103 670
use contact$4  contact$4_0
array 0 9 1000 0 0 0
timestamp 1635942583
transform 1 0 -781 0 1 -1885
box -64 -32 64 32
<< end >>
